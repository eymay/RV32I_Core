module immed_gen_tb ();
    
    

endmodule